module LF1 (input [31:0] data, output [31:0] out);
   
   assign out = data << 1;
   
endmodule 
