module MyAnd
(
   input [31:0]  x,
                 y,
					  
	
   output [31:0] A
);

and and1 [31:0] (A,x,y);

endmodule