module MyOr
(
   input [31:0]  x,
                 y,
					  
	
   output [31:0] A
);

or or1 [31:0] (A,x,y);

endmodule